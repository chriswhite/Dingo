["Fast Cars", "Weightlifting"]  |  {"name": {"first": "Joe", "last": "Sixpack"}, "gender": "MALE", "age": 30, "verified": false}
["Fashion", "Food", "Yoga"]     |  {"name": {"first": "Jane", "last": "Curvey"}, "gender": "FEMALE", "age": 25, "verified": true}