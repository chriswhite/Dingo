0.5	|	4	|	3	|	2	|	1
-7.5	|	5	|	10	|	20	|	30
14	|	20	|	10	|	2.5	|	3.5